library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.numeric_std.all;

entity InstructionMemory is
    Port ( Address : in STD_LOGIC_VECTOR (7 downto 0);
           DataOut : out STD_LOGIC_VECTOR (31 downto 0));
end InstructionMemory;

architecture Structural of InstructionMemory is
type storage_type is array (0 to 63) of std_logic_vector(31 downto 0);

-- COMENTAR A LINHA SEGUINTE E DESCOMENTAR AS LINHAS CORRESPONDENTES AO TURNO DA SEMANA
--signal storage: storage_type := (others => x"00000000");

----------------------------------------------------------------------------------------------------
-- MEMORY
----------------------------------------------------------------------------------------------------
signal storage: storage_type := (
          --    OPCODE &   DR   &   SA   &   SB   &        KNS        -- ASSEMBLY CODE
        -- 0 => "000001" & "0001" & "0000" & "1111" & "11010011000011", --        ADDI  R1,R0,#-2876
         --1 => "000001" & "0111" & "0000" & "1111" & "11111111111000", --        ADDI  R7,R0,#-8
         --2 => "000001" & "0010" & "0000" & "0000" & "00000000001111", --        ADDI  R2,R0,#15
         --3 => "001100" & "0011" & "0000" & "0000" & "00000000000000", --        XOR   R3,R0,R0
         --4 => "001100" & "0100" & "0001" & "0010" & "00000000000000", -- LOOP:  XOR   R4,R1,R2
         --5 => "000100" & "0100" & "0100" & "0010" & "00000000000000", --        AND   R4,R4,R2
         --6 => "010100" & "0101" & "0100" & "0000" & "00000000000000", --        LD    R5,(R4+R0)
         --7 => "010011" & "0001" & "0000" & "0001" & "00000000000000", --        SHRA  R1,R1
         --8 => "010011" & "0001" & "0000" & "0001" & "00000000000000", --        SHRA  R1,R1
         --9 => "010011" & "0001" & "0000" & "0001" & "00000000000000", --        SHRA  R1,R1
        --10 => "010011" & "0001" & "0000" & "0001" & "00000000000000", --        SHRA  R1,R1
        --11 => "000000" & "0011" & "0011" & "0101" & "00000000000000", --        ADD   R3,R3,R5
        --12 => "011000" & "0011" & "0001" & "0111" & "11111111111111", --        BI.NE R1,#-1,R7     ; --> if (R4 >= R3) goto LOOP
        --13 => "010111" & "1001" & "0000" & "0000" & "00000000000000", -- END:   B     #0            ; --> END
           -
           --TESTING PROB
           -- 0=> "00000101010000000000000000001010",
            --1=>"00000101100000000000000000000000",
            --2=>"01011000000110010100000000000000",
            --3=>"00000101010000000000000000010100",
            --4=>"01011000000110010100000000000100",
            --5=>"01010100010110000000000000000000",
            --6=>"01010100100110000000000000000100",
            --7=>"00001000110010000100000000000000",
            --8=>"01011101010011000000000000000010",
            --9=>"00001000110001001000000000000000",
            --10=>"01011000000110001100000000001000",
            --11=>"010111" & "1001" & "0000" & "0000" & "00000000000000",
     0 => "00000100010000000000001000000000",   --  ADDI    R1,R0,#512
     1 => "00000100100000000000000000000001",   --  ADDI    R2,R0,#1
     2 => "01011000000001001000000000000000",   --  ST      0(R1),R2
     3 => "00000000010001001000000000000000",   --  ADD     R1,R1,R2
     4 => "01011000000001001000000000000000",   --  ST      0(R1),R2
     5 => "00001100110001111111111111110110",   --  SUBI    R3,R1,#-10
     6 => "00000111100000000000010000000000",   --  ADDI    R14,R0,#1024
     7 => "01010001000001000000000000000000",   --  LD      R4,R0(R1)
     8 => "01010101010001111111111111111111",   --  LDI     R5,-1(R1)
     9 => "00000001100100010100000000000000",   --  ADD     R6,R4,R5
    10 => "01011000000001011000000000000001",   --  ST      1(R1),R6
    11 => "00000100010001000000000000000001",   --  ADDI    R1,R1,#1
    12 => "01011100110001001111111111111011",   --  B.NEQ   -5,R1,R3
    13 => "00000100110000000000001000000000",   --  ADDI    R3,R0,#512
    14 => "00001010000011000100000000000000",   --  SUB     R8,R3,R1
    15 => "01010101110001000000000000000000",   --  LDI     R7,0(R1)
    16 => "00000111010000000000000000010100",   --  ADDI    R13,R0,#20
    17 => "01101011101000110100000000000000",   --  JIL.LT  R13,R8,0
    18 => "01011100100100010000000000001001",   --  B.EQ    9,R4,R4
    19 => "00000000000000000000000000000000",   --  ADD     R0,R0,R0
    20 => "00000100100010000000000000000001",   --  ADDI    R2,R2,#1
    21 => "01010110010001111111111111111111",   --  LDI     R9,-1(R1)
    22 => "00000001110111100100000000000000",   --  ADD     R7,R7,R9
    23 => "00001100010001000000000000000001",   --  SUBI    R1,R1,#1
    24 => "00000110001000000000000000000001",   --  ADDI    R8,R8,#1
    25 => "00000111111111111111111111111111",   --  ADDI    R15,R15,#-1
    26 => "01101000010000111100000000000000",   --  JI      
    27 => "01011110010000000000000000000001",   --  BL      1
    28 => "01101000010000111100000000000000",   --  JI      R15
   -- others => "00000000000000000000000000000000"   --  NOP

    others => x"00000000" -- NOP
	 );

	 
begin

DataOut <= storage(to_integer(unsigned(Address)));
	
end Structural;
